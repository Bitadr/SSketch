`timescale 1ns / 1ps


module omp_test();

parameter P =  16;

reg 	clk;
reg 	rst;
reg   ap_start;
wire   ap_done;
wire   ap_idle;
wire   ap_ready;

wire  [10:0] Q_address0[P-1:0];
wire   Q_ce0[P-1:0];
wire   Q_we0[P-1:0];
wire  [31:0] Q_d0[P-1:0];
reg [31:0] Q_q0[P-1:0];



/*wire  [14:0] Q_address0[P-1:0];
wire   Q_ce0[P-1:0];
wire   Q_we0[P-1:0];
wire  [31:0] Q_d0[P-1:0];
wire [31:0] Q_q0[P-1:0];*/



wire  [7:0] X_address0;
wire   X_ce0;
reg [31:0] X_q0;
wire [31:0] X_d0;
wire X_we0;


reg  [31:0] l;
reg  [31:0] k;
reg  [31:0] epsilon;

wire  [6:0] V_address0;
wire   V_ce0;
wire   V_we0;
wire  [31:0] V_d0;
wire  [31:0] V_q0;

wire  [6:0] supp_address0;
wire   supp_ce0;
wire   supp_we0;
wire  [31:0] supp_d0;
wire [31:0] supp_q0;

wire  [31:0] supp_len;
wire   supp_len_ap_vld;








/*always @(posedge clk)
	X_q0 <= {X_address0, 14'b0} + 32'h3DCCCCCD;*/

reg  [10:0] Q_address[P-1:0];
reg   Q_we[P-1:0];
reg  [31:0] Q_d[P-1:0];



/*reg  [14:0] Q_address[P-1:0];
reg   Q_we[P-1:0];
reg  [31:0] Q_d[P-1:0];*/





reg g;	
		

omp_supp suppRAM (
  .clka(clk), // input clka
  .wea(supp_we0), // input [0 : 0] wea
  .addra(supp_address0), // input [6 : 0] addra
  .dina(supp_d0), // input [31 : 0] dina
  .douta(supp_q0) // output [31 : 0] douta
);
	

omp_V VRAM (
  .clka(clk), // input clka
  .wea(V_we0), // input [0 : 0] wea
  .addra(V_address0), // input [6 : 0] addra
  .dina(V_d0), // input [31 : 0] dina
  .douta(V_q0) // output [31 : 0] douta
);	



	reg [31:0]Q_mem [P-1:0] [2047:0];
	//reg [31:0] X_mem [255:0];


	
	
//			always @(posedge clk)
//		begin
//			X_q0 <= X_mem[ X_address0];
//		end
		
		


genvar i;
generate
	for(i=0;i<P;i=i+1)
	begin:MEM
//	omp_Q Q_u (
//  .clka(clk), // input clka
//  .wea(g? Q_we[i] : Q_we0[i]), // input [0 : 0] wea
//  .addra(g? Q_address[i]: Q_address0[i]), // input [10 : 0] addra
//  .dina(g? Q_d[i]:Q_d0[i]), // input [31 : 0] dina
//  .douta(Q_q0[i]) // output [31 : 0] douta
//);	

		always @(posedge clk)
		begin
			if(g? Q_we[i] : Q_we0[i])
			begin
					Q_mem[i][ g? Q_address[i]: Q_address0[i]] <= g? 32'b0:Q_d0[i];
			end
			Q_q0[i] <= Q_mem[i][g? Q_address[i]: Q_address0[i]];
		end
	end

endgenerate



integer j,kk;
initial begin
		clk = 0;
		rst = 1;
		ap_start = 0;
		epsilon = 32'h3dcccccd;
		k = 32'd100;
		l = 32'd100;
		g=1;
//	$readmemh("X",X_mem);
	
/*$readmemh("Q0",Q_mem[0]);
$readmemh("Q1",Q_mem[1]);
$readmemh("Q2",Q_mem[2]);
$readmemh("Q3",Q_mem[3]);
$readmemh("Q4",Q_mem[4]);
$readmemh("Q5",Q_mem[5]);
$readmemh("Q6",Q_mem[6]);
$readmemh("Q7",Q_mem[7]);
$readmemh("Q8",Q_mem[8]);
$readmemh("Q9",Q_mem[9]);
$readmemh("Q10",Q_mem[10]);
$readmemh("Q11",Q_mem[11]);
$readmemh("Q12",Q_mem[12]);
$readmemh("Q13",Q_mem[13]);
$readmemh("Q14",Q_mem[14]);
$readmemh("Q15",Q_mem[15]);*/
	

		#1000
		rst = 0;
		g=0;
		@(negedge clk)
		ap_start = 1;
		//@(negedge clk)
	//	ap_start =0;
		@(negedge ap_done);
		#1000
		$finish;
	end

	always #5 clk = ~clk;


omp omp_uut (
    .ap_clk(clk), 
    .ap_rst(rst), 
    .ap_start(ap_start), 
    .ap_done(ap_done), 
    .ap_idle(ap_idle), 
    .ap_ready(ap_ready), 
	
    .Qt_0_address0(Q_address0[0]), 
    .Qt_0_ce0(Q_ce0[0]), 
    .Qt_0_we0(Q_we0[0]), 
    .Qt_0_d0(Q_d0[0]), 
    .Qt_0_q0(Q_q0[0]), 
	
	.Qt_1_address0(Q_address0[1]), 
    .Qt_1_ce0(Q_ce0[1]), 
    .Qt_1_we0(Q_we0[1]), 
    .Qt_1_d0(Q_d0[1]), 
    .Qt_1_q0(Q_q0[1]), 
	
	.Qt_2_address0(Q_address0[2]), 
    .Qt_2_ce0(Q_ce0[2]), 
    .Qt_2_we0(Q_we0[2]), 
    .Qt_2_d0(Q_d0[2]), 
    .Qt_2_q0(Q_q0[2]), 
	
	.Qt_3_address0(Q_address0[3]), 
    .Qt_3_ce0(Q_ce0[3]), 
    .Qt_3_we0(Q_we0[3]), 
    .Qt_3_d0(Q_d0[3]), 
    .Qt_3_q0(Q_q0[3]), 
	
	.Qt_4_address0(Q_address0[4]), 
    .Qt_4_ce0(Q_ce0[4]), 
    .Qt_4_we0(Q_we0[4]), 
    .Qt_4_d0(Q_d0[4]), 
    .Qt_4_q0(Q_q0[4]), 
	
	.Qt_5_address0(Q_address0[5]), 
    .Qt_5_ce0(Q_ce0[5]), 
    .Qt_5_we0(Q_we0[5]), 
    .Qt_5_d0(Q_d0[5]), 
    .Qt_5_q0(Q_q0[5]), 
	
	.Qt_6_address0(Q_address0[6]), 
    .Qt_6_ce0(Q_ce0[6]), 
    .Qt_6_we0(Q_we0[6]), 
    .Qt_6_d0(Q_d0[6]), 
    .Qt_6_q0(Q_q0[6]), 
	
	.Qt_7_address0(Q_address0[7]), 
    .Qt_7_ce0(Q_ce0[7]), 
    .Qt_7_we0(Q_we0[7]), 
    .Qt_7_d0(Q_d0[7]), 
    .Qt_7_q0(Q_q0[7]), 
	
	.Qt_8_address0(Q_address0[8]), 
    .Qt_8_ce0(Q_ce0[8]), 
    .Qt_8_we0(Q_we0[8]), 
    .Qt_8_d0(Q_d0[8]), 
    .Qt_8_q0(Q_q0[8]), 
	
	.Qt_9_address0(Q_address0[9]), 
    .Qt_9_ce0(Q_ce0[9]), 
    .Qt_9_we0(Q_we0[9]), 
    .Qt_9_d0(Q_d0[9]), 
    .Qt_9_q0(Q_q0[9]), 
	
	.Qt_10_address0(Q_address0[10]), 
    .Qt_10_ce0(Q_ce0[10]), 
    .Qt_10_we0(Q_we0[10]), 
    .Qt_10_d0(Q_d0[10]), 
    .Qt_10_q0(Q_q0[10]), 
	
	.Qt_11_address0(Q_address0[11]), 
    .Qt_11_ce0(Q_ce0[11]), 
    .Qt_11_we0(Q_we0[11]), 
    .Qt_11_d0(Q_d0[11]), 
    .Qt_11_q0(Q_q0[11]), 
	
	.Qt_12_address0(Q_address0[12]), 
    .Qt_12_ce0(Q_ce0[12]), 
    .Qt_12_we0(Q_we0[12]), 
    .Qt_12_d0(Q_d0[12]), 
    .Qt_12_q0(Q_q0[12]), 
	
	.Qt_13_address0(Q_address0[13]), 
    .Qt_13_ce0(Q_ce0[13]), 
    .Qt_13_we0(Q_we0[13]), 
    .Qt_13_d0(Q_d0[13]), 
    .Qt_13_q0(Q_q0[13]), 
	
	.Qt_14_address0(Q_address0[14]), 
    .Qt_14_ce0(Q_ce0[14]), 
    .Qt_14_we0(Q_we0[14]), 
    .Qt_14_d0(Q_d0[14]), 
    .Qt_14_q0(Q_q0[14]), 
	
	.Qt_15_address0(Q_address0[15]), 
    .Qt_15_ce0(Q_ce0[15]), 
    .Qt_15_we0(Q_we0[15]), 
    .Qt_15_d0(Q_d0[15]), 
    .Qt_15_q0(Q_q0[15]), 
	
    .X_address0(X_address0), 
    .X_ce0(X_ce0), 
    .X_q0(X_q0), 

    .l(l), 
    .k(k), 
    .epsilon(epsilon), 
    .V_address0(V_address0), 
    .V_ce0(V_ce0), 
    .V_we0(V_we0), 
    .V_d0(V_d0), 
   .V_q0(V_q0), 
    .supp_address0(supp_address0), 
    .supp_ce0(supp_ce0), 
    .supp_we0(supp_we0), 
    .supp_d0(supp_d0), 
    .supp_q0(supp_q0), 
    .supp_len(supp_len),
    .supp_len_ap_vld(supp_len_ap_vld)
    );
	/* omp instance_name (
   
    .ap_clk(clk), 
    .ap_rst(rst), 
    .ap_start(ap_start), 
    .ap_done(ap_done), 
    .ap_idle(ap_idle), 
    .ap_ready(ap_ready), 
	
    .Qt_address0(Q_address0[0]), 
    .Qt_ce0(Q_ce0[0]), 
    .Qt_we0(Q_we0[0]), 
    .Qt_d0(Q_d0[0]), 
    .Qt_q0(Q_q0[0]), 
	 
	 .X_address0(X_address0), 
    .X_ce0(X_ce0), 
    .X_q0(X_q0), 

    .l(l), 
    .k(k), 
    .epsilon(epsilon), 
    .V_address0(V_address0), 
    .V_ce0(V_ce0), 
    .V_we0(V_we0), 
    .V_d0(V_d0), 
    .V_q0(V_q0), 
    .supp_address0(supp_address0), 
    .supp_ce0(supp_ce0), 
    .supp_we0(supp_we0), 
    .supp_d0(supp_d0), 
    .supp_q0(supp_q0), 
    .supp_len(supp_len),
.supp_len_ap_vld(supp_len_ap_vld));*/




 

endmodule
